module storage()

//get written to by camera_interface

//store written data

//get read by hdmi_interface